
// instr_mem.v - instruction memory for single-cycle MIPS32 CPU

module instr_mem #(parameter DATA_WIDTH = 32, ADDR_WIDTH = 6, MEM_SIZE = 64) (
    input       [ADDR_WIDTH-1:0] instr_addr,
    output      [DATA_WIDTH-1:0] instr
);

// array of 64 32-bit words or instructions
reg [DATA_WIDTH-1:0] instr_ram [0:MEM_SIZE-1];

initial begin
    $readmemh("program_dump.hex", instr_ram);
end

// word-aligned memory access
// combinational read logic
assign instr = instr_ram[instr_addr];

endmodule
