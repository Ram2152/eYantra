
// alu.v - ALU module

module alu #(parameter WIDTH = 32) (
    input       [WIDTH-1:0] a, b,       // operands
    input       [2:0] alu_ctrl,         // ALU control
    output reg  [WIDTH-1:0] alu_out,    // ALU output
    output      zero                    // zero flag
);

always @(a, b, alu_ctrl) begin
    case (alu_ctrl)
        3'b000: alu_out <= a & b;         // AND
        3'b001: alu_out <= a | b;         // OR
        3'b010: alu_out <= a + b;         // ADD
        3'b110: alu_out <= a + ~b + 1;    // SUB
        3'b111: if (a[31] != b[31])       // SLT
                    alu_out <= a[31] ? 0 : 1;
                else
                    alu_out <= a < b ? 1 : 0;
        default: alu_out = 0;
    endcase
end

assign zero = (alu_out == 0);

endmodule
